LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

USE work.fLink_definitions.ALL;

PACKAGE mpc5200b_to_axi_master_pkg IS
	CONSTANT c_axi_id_width	: INTEGER := 1;
	CONSTANT c_burst_type_fixed	: STD_LOGIC_VECTOR := "00";
	CONSTANT c_burst_type_incr	: STD_LOGIC_VECTOR := "01";
	CONSTANT c_burst_type_wrap	: STD_LOGIC_VECTOR := "10";
	CONSTANT c_address_width : INTEGER := 32;
	
	COMPONENT lpb_mpc5200b_to_axi_master IS
		GENERIC (
			LPBADDRWIDTH 	: INTEGER := 32;
			LPBDATAWIDTH	: INTEGER := 32;
			LPBTSIZEWIDTH	: INTEGER := 3;
			LPBCSWIDTH		: INTEGER := 2;
			LPBBANKWIDTH	: INTEGER := 2
		);
		PORT (
			-- Clock and Reset
			clk			:   IN  STD_LOGIC;
			reset_n		: 	IN  STD_LOGIC;

			-- Write Address Channel
			axi_awid 			: OUT STD_LOGIC_VECTOR(c_axi_id_width-1 downto 0); -- Write Address ID
			axi_awaddr 			: OUT STD_LOGIC_VECTOR(c_address_width-1 downto 0); -- Write address
			axi_awlen 			: OUT STD_LOGIC_VECTOR(7 downto 0); -- Burst length. The burst length gives the exact number of transfers in a burst
			axi_awsize 			: OUT STD_LOGIC_VECTOR(2 downto 0); -- Burst size. This signal indicates the size of each transfer in the burst
			axi_awburst 		: OUT STD_LOGIC_VECTOR(1 downto 0); -- Burst type. The burst type and the size information, determine how the address for each transfer within the burst is calculated.
			axi_awvalid 		: OUT STD_LOGIC; -- Write address valid. This signal indicates that the channel is signaling valid write address and control information.
			axi_awready 		: IN STD_LOGIC; -- Write address ready. This signal indicates that the slave is ready to accept an address and associated control signals.
			axi_awprot 			: OUT STD_LOGIC_VECTOR(2 downto 0); --Protection type. This signal indicates the privilege and security level of the transaction, and whether the transaction is a data access or an instruction access.

			-- Write Data Channel
			axi_wdata 			: OUT STD_LOGIC_VECTOR(c_fLink_avs_data_width-1 downto 0); -- Write Data
			axi_wstrb 			: OUT STD_LOGIC_VECTOR(3 downto 0); -- Write strobes. This signal indicates which byte lanes hold valid data. There is one write strobe bit for each eight bits of the write data bus.
			axi_wvalid 			: OUT STD_LOGIC; -- Write valid. This signal indicates that valid write data and strobes are available.
			axi_wready 			: IN STD_LOGIC; -- Write ready. This signal indicates that the slave can accept the write data.
			axi_wlast			: OUT STD_LOGIC; --Write last. This signal indicates the last transfer in a write burst
			
			
			-- Read Address Channel
			axi_araddr 			: OUT STD_LOGIC_VECTOR(c_address_width-1 downto 0); -- Read address. This signal indicates the initial address of a read burst transaction.
			axi_arvalid 		: OUT STD_LOGIC; -- Read address valid. This signal indicates that the channel is signaling valid read address and control information.
			axi_arready			: IN STD_LOGIC; -- Read address ready. This signal indicates that the slave is ready to accept an address and associated  control signals.
			axi_arid 			: OUT STD_LOGIC_VECTOR(c_axi_id_width-1 downto 0); -- Read address ID. This signal is the identification tag for the read address group of signals.
			axi_arlen 			: OUT STD_LOGIC_VECTOR(7 downto 0); -- Burst length. The burst length gives the exact number of transfers in a burst
			axi_arsize 			: OUT STD_LOGIC_VECTOR(2 downto 0); -- Burst size. This signal indicates the size of each transfer in the burst
			axi_arburst 		: OUT STD_LOGIC_VECTOR(1 downto 0); -- Burst type. The burst type and the size information,  determine how the address for each transfer within the burst is calculated.
			axi_arprot 			: OUT STD_LOGIC_VECTOR(2 downto 0); --Protection type. This signal indicates the privilege and security level of the transaction, and whether the transaction is a data access or an instruction access
			-- Read Data Channel
			axi_rdata 			: IN STD_LOGIC_VECTOR(c_fLink_avs_data_width-1 downto 0); -- Read Data
			axi_rresp 			: IN STD_LOGIC_VECTOR(1 downto 0); -- Read response. This signal indicates the status of the read transfer.
			axi_rvalid 			: IN STD_LOGIC; -- Read valid. This signal indicates that the channel is signaling the required read data.
			axi_rready 			: OUT STD_LOGIC; -- Read ready. This signal indicates that the master can accept the read data and response information
			axi_rid 			: IN STD_LOGIC_VECTOR(c_axi_id_width-1 downto 0); -- Read ID tag. This signal is the identification tag for the read data group of signals generated by the slave.
			axi_rlast 			: IN STD_LOGIC; -- Read last. This signal indicates the last transfer in a read burst.
			-- Write Response Channel
			axi_bresp 			: IN STD_LOGIC_VECTOR(1 downto 0); -- Write response. This signal indicates the status of the write transaction.
			axi_bvalid 			: IN STD_LOGIC; -- Write response valid. This signal indicates that the channel is signaling a valid write response.
			axi_bready 			: OUT STD_LOGIC;	-- Response ready. This signal indicates that the master can accept a write response.
			axi_bid 			: IN STD_LOGIC_VECTOR(c_axi_id_width-1 downto 0); -- Response ID tag. This signal is the ID tag of the write response.
			
			-- LocalPlus signals
			lpb_ad		: 	INOUT	STD_LOGIC_VECTOR ((LPBDATAWIDTH-1) DOWNTO 0);
			lpb_cs_n	: 	IN	STD_LOGIC_VECTOR ((LPBCSWIDTH-1) DOWNTO 0);
			lpb_oe_n	: 	IN	STD_LOGIC;
			lpb_ack_n	: 	OUT	STD_LOGIC;
			lpb_ale_n	: 	IN	STD_LOGIC;
			lpb_rdwr_n	: 	IN	STD_LOGIC;
			lpb_ts_n	: 	IN	STD_LOGIC
		);
	END COMPONENT;	

END PACKAGE mpc5200b_to_axi_master_pkg;



LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
USE work.mpc5200b_to_axi_master_pkg.ALL;
USE work.fLink_definitions.ALL;

ENTITY lpb_mpc5200b_to_axi_master IS
	
	GENERIC (
			LPBADDRWIDTH 	: INTEGER := 32;
			LPBDATAWIDTH	: INTEGER := 32;
			LPBTSIZEWIDTH	: INTEGER := 3;
			LPBCSWIDTH		: INTEGER := 2;
			LPBBANKWIDTH	: INTEGER := 2
		);
		PORT (
			-- Clock and Reset
			clk			:   IN  STD_LOGIC;
			reset_n		: 	IN  STD_LOGIC;

			-- Write Address Channel
			axi_awid 			: OUT STD_LOGIC_VECTOR(c_axi_id_width-1 downto 0); -- Write Address ID
			axi_awaddr 			: OUT STD_LOGIC_VECTOR(c_address_width-1 downto 0); -- Write address
			axi_awlen 			: OUT STD_LOGIC_VECTOR(7 downto 0); -- Burst length. The burst length gives the exact number of transfers in a burst
			axi_awsize 			: OUT STD_LOGIC_VECTOR(2 downto 0); -- Burst size. This signal indicates the size of each transfer in the burst
			axi_awburst 		: OUT STD_LOGIC_VECTOR(1 downto 0); -- Burst type. The burst type and the size information, determine how the address for each transfer within the burst is calculated.
			axi_awvalid 		: OUT STD_LOGIC; -- Write address valid. This signal indicates that the channel is signaling valid write address and control information.
			axi_awready 		: IN STD_LOGIC; -- Write address ready. This signal indicates that the slave is ready to accept an address and associated control signals.
			axi_awprot 			: OUT STD_LOGIC_VECTOR(2 downto 0); --Protection type. This signal indicates the privilege and security level of the transaction, and whether the transaction is a data access or an instruction access.

			-- Write Data Channel
			axi_wdata 			: OUT STD_LOGIC_VECTOR(c_fLink_avs_data_width-1 downto 0); -- Write Data
			axi_wstrb 			: OUT STD_LOGIC_VECTOR(3 downto 0); -- Write strobes. This signal indicates which byte lanes hold valid data. There is one write strobe bit for each eight bits of the write data bus.
			axi_wvalid 			: OUT STD_LOGIC; -- Write valid. This signal indicates that valid write data and strobes are available.
			axi_wready 			: IN STD_LOGIC; -- Write ready. This signal indicates that the slave can accept the write data.
			axi_wlast			: OUT STD_LOGIC; --Write last. This signal indicates the last transfer in a write burst
			
			
			-- Read Address Channel
			axi_araddr 			: OUT STD_LOGIC_VECTOR(c_address_width-1 downto 0); -- Read address. This signal indicates the initial address of a read burst transaction.
			axi_arvalid 		: OUT STD_LOGIC; -- Read address valid. This signal indicates that the channel is signaling valid read address and control information.
			axi_arready			: IN STD_LOGIC; -- Read address ready. This signal indicates that the slave is ready to accept an address and associated  control signals.
			axi_arid 			: OUT STD_LOGIC_VECTOR(c_axi_id_width-1 downto 0); -- Read address ID. This signal is the identification tag for the read address group of signals.
			axi_arlen 			: OUT STD_LOGIC_VECTOR(7 downto 0); -- Burst length. The burst length gives the exact number of transfers in a burst
			axi_arsize 			: OUT STD_LOGIC_VECTOR(2 downto 0); -- Burst size. This signal indicates the size of each transfer in the burst
			axi_arburst 		: OUT STD_LOGIC_VECTOR(1 downto 0); -- Burst type. The burst type and the size information,  determine how the address for each transfer within the burst is calculated.
			axi_arprot 			: OUT STD_LOGIC_VECTOR(2 downto 0); --Protection type. This signal indicates the privilege and security level of the transaction, and whether the transaction is a data access or an instruction access
			-- Read Data Channel
			axi_rdata 			: IN STD_LOGIC_VECTOR(c_fLink_avs_data_width-1 downto 0); -- Read Data
			axi_rresp 			: IN STD_LOGIC_VECTOR(1 downto 0); -- Read response. This signal indicates the status of the read transfer.
			axi_rvalid 			: IN STD_LOGIC; -- Read valid. This signal indicates that the channel is signaling the required read data.
			axi_rready 			: OUT STD_LOGIC; -- Read ready. This signal indicates that the master can accept the read data and response information
			axi_rid 			: IN STD_LOGIC_VECTOR(c_axi_id_width-1 downto 0); -- Read ID tag. This signal is the identification tag for the read data group of signals generated by the slave.
			axi_rlast 			: IN STD_LOGIC; -- Read last. This signal indicates the last transfer in a read burst.
			-- Write Response Channel
			axi_bresp 			: IN STD_LOGIC_VECTOR(1 downto 0); -- Write response. This signal indicates the status of the write transaction.
			axi_bvalid 			: IN STD_LOGIC; -- Write response valid. This signal indicates that the channel is signaling a valid write response.
			axi_bready 			: OUT STD_LOGIC;	-- Response ready. This signal indicates that the master can accept a write response.
			axi_bid 			: IN STD_LOGIC_VECTOR(c_axi_id_width-1 downto 0); -- Response ID tag. This signal is the ID tag of the write response.
			
			-- LocalPlus signals
			lpb_ad		: 	INOUT	STD_LOGIC_VECTOR ((LPBDATAWIDTH-1) DOWNTO 0);
			lpb_cs_n	: 	IN	STD_LOGIC_VECTOR ((LPBCSWIDTH-1) DOWNTO 0);
			lpb_oe_n	: 	IN	STD_LOGIC;
			lpb_ack_n	: 	OUT	STD_LOGIC;
			lpb_ale_n	: 	IN	STD_LOGIC;
			lpb_rdwr_n	: 	IN	STD_LOGIC;
			lpb_ts_n	: 	IN	STD_LOGIC
		);
END lpb_mpc5200b_to_axi_master;

---------------------------------------------------------

-- reset SIGNAL einbauen

---------------------------------------------------------

ARCHITECTURE rtl OF lpb_mpc5200b_to_axi_master IS

SIGNAL lpb_adr_q 			: STD_LOGIC_VECTOR((LPBADDRWIDTH-1) DOWNTO 0);
SIGNAL lpb_data_q			: STD_LOGIC_VECTOR((LPBDATAWIDTH-1) DOWNTO 0);
SIGNAL lpb_tsize_q 			: STD_LOGIC_VECTOR ((LPBTSIZEWIDTH-1) DOWNTO 0);

SIGNAL lpb_data_en			: STD_LOGIC;
SIGNAL lpb_start			: STD_LOGIC;

SIGNAL lpb_rd				: STD_LOGIC;
SIGNAL lpb_wr				: STD_LOGIC;
SIGNAL lpb_ack_i			: STD_LOGIC;

SIGNAL lpb_start_en			: STD_LOGIC;

SIGNAL lpb_ad_o				: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL lpb_ad_en			: STD_LOGIC;

SIGNAL arvalid_i			: STD_LOGIC := '0';
SIGNAL awvalid_i			: STD_LOGIC := '0';

type state IS (init, act, rst);
SIGNAL axistate 			: state;

BEGIN
--activation of FPGA with only one chip select SIGNAL
lpb_rd <= (NOT lpb_cs_n(0) AND NOT lpb_oe_n);
lpb_wr <= (NOT lpb_cs_n(0) AND NOT lpb_rdwr_n);

-- external ack SIGNAL gets internal value
lpb_ack_n <= NOT lpb_ack_i;

axi_awid <= (OTHERS =>'1');
axi_arid <= (OTHERS =>'1');
axi_awprot <= (OTHERS =>'0');
axi_arprot <= (OTHERS =>'0');
-- ############################# MPC interface functions ##############################
-- tristate buffer generation

lpb_data_switching : PROCESS(lpb_ad_o, lpb_ad_en, reset_n)
	BEGIN
		IF reset_n = '0' THEN
			lpb_ad <= (OTHERS => 'Z');
		ELSIF lpb_ad_en = '1' THEN
				lpb_ad <= lpb_ad_o;
		ELSE
				lpb_ad <= (OTHERS => 'Z');
		END IF;
	END PROCESS;


-- mpc_address_latching : necessary because of multiplexed bus system
-- latching of addresses at falling edge of clk

lpb_address_latching : PROCESS (clk, reset_n)

	BEGIN
		IF reset_n = '0' THEN
			lpb_adr_q <= (OTHERS => '0');
			lpb_tsize_q <= (OTHERS => '0');
		ELSIF rising_edge(clk) THEN									
			IF lpb_ale_n = '0' THEN
				lpb_adr_q <= lpb_ad((LPBADDRWIDTH-1) DOWNTO 0);
				lpb_tsize_q   <= lpb_ad((LPBDATAWIDTH-2) DOWNTO (LPBDATAWIDTH-4));
			END IF;	
		END IF;	
		
	END PROCESS lpb_address_latching;

-- lpb_write_data_latching
-- latching of data of the lpb bus at write cycle

lpb_write_data_latching : PROCESS (clk, reset_n)			

	BEGIN
		IF reset_n = '0' THEN
			lpb_data_q <= (OTHERS => '0');
			lpb_data_en <= '0';
			lpb_start <= '0';
		ELSE
			IF rising_edge (clk) THEN
				IF lpb_ts_n = '0' AND lpb_start = '0' THEN
					--lpb_start <= '1';		-- for 66MHz we can start here
					lpb_start_en <= '1';
				ELSE
					--lpb_start <= '0';
					lpb_start_en <= '0';
				END IF;
				
				-- needable for 33MHz support, for 66MHz we can start erlier
				IF lpb_start_en = '1' THEN
					lpb_start <= '1';
				ELSE	
					lpb_start <= '0';
				END IF;
					
				IF lpb_ts_n = '0' AND lpb_rdwr_n = '0' THEN
					lpb_data_en <= '1';				-- wait 1 clock cycle for data ready
				END IF;
			
				IF lpb_data_en = '1' THEN
					lpb_data_q <= lpb_ad;
					lpb_data_en <= '0';				
				END IF;
			END IF;
		END IF;
END PROCESS lpb_write_data_latching;

axi_read_address_channel : PROCESS (reset_n, clk)
	BEGIN
		IF reset_n = '0' THEN
			axi_arvalid <= '0';
			arvalid_i <= '0';
			axi_araddr <= (OTHERS => '0');
			axi_arlen 	<= "00000000";	--only one transfer
			axi_arsize 	<= "010";
			axi_arburst <= "01"; --increment	
		ELSIF rising_edge(clk) THEN	
			IF lpb_start = '1' AND lpb_rd = '1' THEN --start read transfer
				axi_araddr <= lpb_adr_q;
				axi_arvalid <= '1';		
				arvalid_i <= '1';				
			ELSIF(arvalid_i = '1' AND axi_arready = '1') THEN
				axi_arvalid <= '0';
				arvalid_i <= '0';
				axi_araddr <= (OTHERS => '0');
			END IF;
		END IF;
END PROCESS axi_read_address_channel;

axi_read_data_channel : PROCESS (reset_n, clk)
	BEGIN
		IF reset_n = '0' THEN
			axi_rready <= '0';
			lpb_ad_o <= (OTHERS => '0');
			lpb_ad_en <= '0';
			lpb_ack_i <= '0';	
		ELSIF rising_edge(clk) THEN	
			axi_rready <= '1';
			IF axi_rvalid = '1' THEN --start read transfer
				IF lpb_rd = '1' AND lpb_ack_i = '0' THEN
					lpb_ad_en <= '1';
					lpb_ack_i <= '1';
					lpb_ad_o <=axi_rdata;	
					axi_rready <= '0';
				END IF;
				
			ELSE
				lpb_ack_i <= '0';	
				lpb_ad_en <= '0';
			END IF;
		END IF;
END PROCESS axi_read_data_channel;

axi_write_address_channel : PROCESS (reset_n, clk)
	BEGIN
		IF reset_n = '0' THEN
			axi_awaddr <= (OTHERS => '0');
			axi_awlen 	<= "00000000";	--only one transfer
			axi_awsize 	<= "010";
			axi_awburst <= "01";
			axi_awvalid <= '0';
		ELSIF rising_edge(clk) THEN	
			IF lpb_start = '1' AND lpb_wr = '1' THEN --start read transfer
				axi_awaddr <= lpb_adr_q;
				axi_awvalid <= '1';		
				awvalid_i <= '1';				
			ELSIF(awvalid_i = '1' AND axi_awready = '1') THEN
				axi_awvalid <= '0';
				awvalid_i <= '0';
				axi_awaddr <= (OTHERS => '0');
			END IF;
		END IF;
END PROCESS axi_write_address_channel;

axi_write_data_channel : PROCESS (reset_n, clk)
	BEGIN
		IF reset_n = '0' THEN
			axi_wstrb <= (OTHERS => '1');
			axi_wdata <= (OTHERS => '0');
			axi_wvalid <= '0';
			axi_wlast <= '0';
		ELSIF rising_edge(clk) THEN	
			IF axi_wready = '1' THEN
				axi_wvalid <= '0';
				axi_wlast <= '0';
			ELSE
				axi_wvalid <= '1';
				axi_wlast <= '1';
				axi_wdata <= lpb_data_q;
			END IF;
		
		END IF;
END PROCESS axi_write_data_channel;

axi_write_response_channel : PROCESS (reset_n, clk)
	BEGIN
		IF reset_n = '0' THEN
			axi_bready <= '1';
		ELSIF rising_edge(clk) THEN	
			IF axi_bvalid = '1' THEN
				axi_bready <= '0';
			ELSE
				axi_bready <= '1';
			END IF;
		END IF;
END PROCESS axi_write_response_channel;

END rtl;